module leftLogicalShiftSixteen(in0, out);
	
	input [31:0] in0;
	output [31:0] out;
	
	assign out[0] = 1'b0;
	assign out[1] = 1'b0;
	assign out[2] = 1'b0;
	assign out[3] = 1'b0;
	assign out[4] = 1'b0;
	assign out[5] = 1'b0;
	assign out[6] = 1'b0;
	assign out[7] = 1'b0;
	assign out[8] = 1'b0;
	assign out[9] = 1'b0;
	assign out[10] = 1'b0;
	assign out[11] = 1'b0;
	assign out[12] = 1'b0;
	assign out[13] = 1'b0;
	assign out[14] = 1'b0;
	assign out[15] = 1'b0;
	assign out[16] = in0[0];
	assign out[17] = in0[1];
	assign out[18] = in0[2];
	assign out[19] = in0[3];
	assign out[20] = in0[4];
	assign out[21] = in0[5];
	assign out[22] = in0[6];
	assign out[23] = in0[7];
	assign out[24] = in0[8];
	assign out[25] = in0[9];
	assign out[26] = in0[10];
	assign out[27] = in0[11];
	assign out[28] = in0[12];
	assign out[29] = in0[13];
	assign out[30] = in0[14];
	assign out[31] = in0[15];

endmodule