module alu_not_33(in0, out);
	
	input [32:0] in0;
	output [32:0] out;
	
	not not_0(out[0], in0[0]);
	not not_1(out[1], in0[1]);
	not not_2(out[2], in0[2]);
	not not_3(out[3], in0[3]);
	not not_4(out[4], in0[4]);
	not not_5(out[5], in0[5]);
	not not_6(out[6], in0[6]);
	not not_7(out[7], in0[7]);
	not not_8(out[8], in0[8]);
	not not_9(out[9], in0[9]);
	not not_10(out[10], in0[10]);
	not not_11(out[11], in0[11]);
	not not_12(out[12], in0[12]);
	not not_13(out[13], in0[13]);
	not not_14(out[14], in0[14]);
	not not_15(out[15], in0[15]);
	not not_16(out[16], in0[16]);
	not not_17(out[17], in0[17]);
	not not_18(out[18], in0[18]);
	not not_19(out[19], in0[19]);
	not not_20(out[20], in0[20]);
	not not_21(out[21], in0[21]);
	not not_22(out[22], in0[22]);
	not not_23(out[23], in0[23]);
	not not_24(out[24], in0[24]);
	not not_25(out[25], in0[25]);
	not not_26(out[26], in0[26]);
	not not_27(out[27], in0[27]);
	not not_28(out[28], in0[28]);
	not not_29(out[29], in0[29]);
	not not_30(out[30], in0[30]);
	not not_31(out[31], in0[31]);
    not not_32(out[32], in0[32]);
	
endmodule
