module rightArithmeticShiftTwo65bit(in0, out);

	input [64:0] in0;
	output [64:0] out;

	assign out[0] = in0[2];
	assign out[1] = in0[3];
	assign out[2] = in0[4];
	assign out[3] = in0[5];
	assign out[4] = in0[6];
	assign out[5] = in0[7];
	assign out[6] = in0[8];
	assign out[7] = in0[9];
	assign out[8] = in0[10];
	assign out[9] = in0[11];
	assign out[10] = in0[12];
	assign out[11] = in0[13];
	assign out[12] = in0[14];
	assign out[13] = in0[15];
	assign out[14] = in0[16];
	assign out[15] = in0[17];
	assign out[16] = in0[18];
	assign out[17] = in0[19];
	assign out[18] = in0[20];
	assign out[19] = in0[21];
	assign out[20] = in0[22];
	assign out[21] = in0[23];
	assign out[22] = in0[24];
	assign out[23] = in0[25];
	assign out[24] = in0[26];
	assign out[25] = in0[27];
	assign out[26] = in0[28];
	assign out[27] = in0[29];
	assign out[28] = in0[30];
	assign out[29] = in0[31];
	assign out[30] = in0[32];
	assign out[31] = in0[33];
	assign out[32] = in0[34];
	assign out[33] = in0[35];
	assign out[34] = in0[36];
	assign out[35] = in0[37];
	assign out[36] = in0[38];
	assign out[37] = in0[39];
	assign out[38] = in0[40];
	assign out[39] = in0[41];
	assign out[40] = in0[42];
	assign out[41] = in0[43];
	assign out[42] = in0[44];
	assign out[43] = in0[45];
	assign out[44] = in0[46];
	assign out[45] = in0[47];
	assign out[46] = in0[48];
	assign out[47] = in0[49];
	assign out[48] = in0[50];
	assign out[49] = in0[51];
	assign out[50] = in0[52];
	assign out[51] = in0[53];
	assign out[52] = in0[54];
	assign out[53] = in0[55];
	assign out[54] = in0[56];
	assign out[55] = in0[57];
	assign out[56] = in0[58];
	assign out[57] = in0[59];
	assign out[58] = in0[60];
	assign out[59] = in0[61];
	assign out[60] = in0[62];
	assign out[61] = in0[63];
	assign out[62] = in0[64];

	assign out[63] = in0[64];
	assign out[64] = in0[64];

endmodule