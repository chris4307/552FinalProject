module register_65(clock, ctrl_writeEnable, ctrl_writeReg, ctrl_readReg, reset, data, out);
	
	input clock, ctrl_writeEnable, reset, ctrl_writeReg, ctrl_readReg;
	input [64:0] data;
	output [64:0] out;


	wire enable_and_reg;
	wire clkn;
	not my_clc_n(clkn, clock);
	//assign enable_and_reg = ctrl_writeReg;
	and my_write_enable_reg_0(enable_and_reg, ctrl_writeEnable, ctrl_writeReg, clkn);

	//module DFFtri(d, clk, clr, pr, in_enable, out_enable, out);
	DFFtri my_dffe_0(.d(data[0]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[0]));
	DFFtri my_dffe_1(.d(data[1]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[1]));
	DFFtri my_dffe_2(.d(data[2]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[2]));
	DFFtri my_dffe_3(.d(data[3]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[3]));
	DFFtri my_dffe_4(.d(data[4]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[4]));
	DFFtri my_dffe_5(.d(data[5]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[5]));
	DFFtri my_dffe_6(.d(data[6]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[6]));
	DFFtri my_dffe_7(.d(data[7]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[7]));
	DFFtri my_dffe_8(.d(data[8]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[8]));
	DFFtri my_dffe_9(.d(data[9]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[9]));
	DFFtri my_dffe_10(.d(data[10]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[10]));
	DFFtri my_dffe_11(.d(data[11]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[11]));
	DFFtri my_dffe_12(.d(data[12]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[12]));
	DFFtri my_dffe_13(.d(data[13]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[13]));
	DFFtri my_dffe_14(.d(data[14]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[14]));
	DFFtri my_dffe_15(.d(data[15]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[15]));
	DFFtri my_dffe_16(.d(data[16]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[16]));
	DFFtri my_dffe_17(.d(data[17]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[17]));
	DFFtri my_dffe_18(.d(data[18]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[18]));
	DFFtri my_dffe_19(.d(data[19]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[19]));
	DFFtri my_dffe_20(.d(data[20]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[20]));
	DFFtri my_dffe_21(.d(data[21]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[21]));
	DFFtri my_dffe_22(.d(data[22]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[22]));
	DFFtri my_dffe_23(.d(data[23]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[23]));
	DFFtri my_dffe_24(.d(data[24]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[24]));
	DFFtri my_dffe_25(.d(data[25]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[25]));
	DFFtri my_dffe_26(.d(data[26]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[26]));
	DFFtri my_dffe_27(.d(data[27]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[27]));
	DFFtri my_dffe_28(.d(data[28]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[28]));
	DFFtri my_dffe_29(.d(data[29]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[29]));
	DFFtri my_dffe_30(.d(data[30]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[30]));
	DFFtri my_dffe_31(.d(data[31]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[31]));
    DFFtri my_dffe_32(.d(data[32]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[32]));
    DFFtri my_dffe_33(.d(data[33]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[33]));
    DFFtri my_dffe_34(.d(data[34]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[34]));
    DFFtri my_dffe_35(.d(data[35]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[35]));
    DFFtri my_dffe_36(.d(data[36]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[36]));
   	DFFtri my_dffe_37(.d(data[37]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[37]));
  	DFFtri my_dffe_38(.d(data[38]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[38]));
	DFFtri my_dffe_39(.d(data[39]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[39]));
	DFFtri my_dffe_40(.d(data[40]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[40]));
	DFFtri my_dffe_41(.d(data[41]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[41]));
	DFFtri my_dffe_42(.d(data[42]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[42]));
	DFFtri my_dffe_43(.d(data[43]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[43]));
	DFFtri my_dffe_44(.d(data[44]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[44]));
	DFFtri my_dffe_45(.d(data[45]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[45]));
	DFFtri my_dffe_46(.d(data[46]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[46]));
	DFFtri my_dffe_47(.d(data[47]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[47]));
	DFFtri my_dffe_48(.d(data[48]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[48]));
	DFFtri my_dffe_49(.d(data[49]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[49]));
	DFFtri my_dffe_50(.d(data[50]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[50]));
	DFFtri my_dffe_51(.d(data[51]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[51]));
	DFFtri my_dffe_52(.d(data[52]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[52]));
	DFFtri my_dffe_53(.d(data[53]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[53]));
	DFFtri my_dffe_54(.d(data[54]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[54]));
	DFFtri my_dffe_55(.d(data[55]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[55]));
	DFFtri my_dffe_56(.d(data[56]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[56]));
	DFFtri my_dffe_57(.d(data[57]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[57]));
	DFFtri my_dffe_58(.d(data[58]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[58]));
	DFFtri my_dffe_59(.d(data[59]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[59]));
	DFFtri my_dffe_60(.d(data[60]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[60]));
	DFFtri my_dffe_61(.d(data[61]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[61]));
	DFFtri my_dffe_62(.d(data[62]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[62]));
	DFFtri my_dffe_63(.d(data[63]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[63]));
	DFFtri my_dffe_64(.d(data[64]), .clk(clock), .clr(reset), .in_enable(enable_and_reg), .out_enable(ctrl_readReg), .out(out[64]));


endmodule
